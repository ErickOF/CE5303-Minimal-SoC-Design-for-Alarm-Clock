// system.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module system (
		output wire       alarm_export,         //         alarm.export
		input  wire       btn_down_export,      //      btn_down.export
		input  wire       btn_set_alarm_export, // btn_set_alarm.export
		input  wire       btn_set_clock_export, // btn_set_clock.export
		input  wire       btn_up_export,        //        btn_up.export
		input  wire       clk_clk,              //           clk.clk
		output wire [3:0] display_h0_export,    //    display_h0.export
		output wire [3:0] display_h1_export,    //    display_h1.export
		output wire [3:0] display_m0_export,    //    display_m0.export
		output wire [3:0] display_m1_export,    //    display_m1.export
		output wire [3:0] display_s0_export,    //    display_s0.export
		output wire [3:0] display_s1_export,    //    display_s1.export
		input  wire       reset_reset_n         //         reset.reset_n
	);

	wire  [31:0] cpu_data_master_readdata;                             // mm_interconnect_0:CPU_data_master_readdata -> CPU:d_readdata
	wire         cpu_data_master_waitrequest;                          // mm_interconnect_0:CPU_data_master_waitrequest -> CPU:d_waitrequest
	wire         cpu_data_master_debugaccess;                          // CPU:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:CPU_data_master_debugaccess
	wire  [14:0] cpu_data_master_address;                              // CPU:d_address -> mm_interconnect_0:CPU_data_master_address
	wire   [3:0] cpu_data_master_byteenable;                           // CPU:d_byteenable -> mm_interconnect_0:CPU_data_master_byteenable
	wire         cpu_data_master_read;                                 // CPU:d_read -> mm_interconnect_0:CPU_data_master_read
	wire         cpu_data_master_write;                                // CPU:d_write -> mm_interconnect_0:CPU_data_master_write
	wire  [31:0] cpu_data_master_writedata;                            // CPU:d_writedata -> mm_interconnect_0:CPU_data_master_writedata
	wire  [31:0] cpu_instruction_master_readdata;                      // mm_interconnect_0:CPU_instruction_master_readdata -> CPU:i_readdata
	wire         cpu_instruction_master_waitrequest;                   // mm_interconnect_0:CPU_instruction_master_waitrequest -> CPU:i_waitrequest
	wire  [14:0] cpu_instruction_master_address;                       // CPU:i_address -> mm_interconnect_0:CPU_instruction_master_address
	wire         cpu_instruction_master_read;                          // CPU:i_read -> mm_interconnect_0:CPU_instruction_master_read
	wire         mm_interconnect_0_uart_avalon_jtag_slave_chipselect;  // mm_interconnect_0:UART_avalon_jtag_slave_chipselect -> UART:av_chipselect
	wire  [31:0] mm_interconnect_0_uart_avalon_jtag_slave_readdata;    // UART:av_readdata -> mm_interconnect_0:UART_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_uart_avalon_jtag_slave_waitrequest; // UART:av_waitrequest -> mm_interconnect_0:UART_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_uart_avalon_jtag_slave_address;     // mm_interconnect_0:UART_avalon_jtag_slave_address -> UART:av_address
	wire         mm_interconnect_0_uart_avalon_jtag_slave_read;        // mm_interconnect_0:UART_avalon_jtag_slave_read -> UART:av_read_n
	wire         mm_interconnect_0_uart_avalon_jtag_slave_write;       // mm_interconnect_0:UART_avalon_jtag_slave_write -> UART:av_write_n
	wire  [31:0] mm_interconnect_0_uart_avalon_jtag_slave_writedata;   // mm_interconnect_0:UART_avalon_jtag_slave_writedata -> UART:av_writedata
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_readdata;       // CPU:debug_mem_slave_readdata -> mm_interconnect_0:CPU_debug_mem_slave_readdata
	wire         mm_interconnect_0_cpu_debug_mem_slave_waitrequest;    // CPU:debug_mem_slave_waitrequest -> mm_interconnect_0:CPU_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_cpu_debug_mem_slave_debugaccess;    // mm_interconnect_0:CPU_debug_mem_slave_debugaccess -> CPU:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_cpu_debug_mem_slave_address;        // mm_interconnect_0:CPU_debug_mem_slave_address -> CPU:debug_mem_slave_address
	wire         mm_interconnect_0_cpu_debug_mem_slave_read;           // mm_interconnect_0:CPU_debug_mem_slave_read -> CPU:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_cpu_debug_mem_slave_byteenable;     // mm_interconnect_0:CPU_debug_mem_slave_byteenable -> CPU:debug_mem_slave_byteenable
	wire         mm_interconnect_0_cpu_debug_mem_slave_write;          // mm_interconnect_0:CPU_debug_mem_slave_write -> CPU:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_writedata;      // mm_interconnect_0:CPU_debug_mem_slave_writedata -> CPU:debug_mem_slave_writedata
	wire         mm_interconnect_0_ram_s1_chipselect;                  // mm_interconnect_0:RAM_s1_chipselect -> RAM:chipselect
	wire  [31:0] mm_interconnect_0_ram_s1_readdata;                    // RAM:readdata -> mm_interconnect_0:RAM_s1_readdata
	wire   [9:0] mm_interconnect_0_ram_s1_address;                     // mm_interconnect_0:RAM_s1_address -> RAM:address
	wire   [3:0] mm_interconnect_0_ram_s1_byteenable;                  // mm_interconnect_0:RAM_s1_byteenable -> RAM:byteenable
	wire         mm_interconnect_0_ram_s1_write;                       // mm_interconnect_0:RAM_s1_write -> RAM:write
	wire  [31:0] mm_interconnect_0_ram_s1_writedata;                   // mm_interconnect_0:RAM_s1_writedata -> RAM:writedata
	wire         mm_interconnect_0_ram_s1_clken;                       // mm_interconnect_0:RAM_s1_clken -> RAM:clken
	wire         mm_interconnect_0_h1_s1_chipselect;                   // mm_interconnect_0:H1_s1_chipselect -> H1:chipselect
	wire  [31:0] mm_interconnect_0_h1_s1_readdata;                     // H1:readdata -> mm_interconnect_0:H1_s1_readdata
	wire   [1:0] mm_interconnect_0_h1_s1_address;                      // mm_interconnect_0:H1_s1_address -> H1:address
	wire         mm_interconnect_0_h1_s1_write;                        // mm_interconnect_0:H1_s1_write -> H1:write_n
	wire  [31:0] mm_interconnect_0_h1_s1_writedata;                    // mm_interconnect_0:H1_s1_writedata -> H1:writedata
	wire         mm_interconnect_0_h0_s1_chipselect;                   // mm_interconnect_0:H0_s1_chipselect -> H0:chipselect
	wire  [31:0] mm_interconnect_0_h0_s1_readdata;                     // H0:readdata -> mm_interconnect_0:H0_s1_readdata
	wire   [1:0] mm_interconnect_0_h0_s1_address;                      // mm_interconnect_0:H0_s1_address -> H0:address
	wire         mm_interconnect_0_h0_s1_write;                        // mm_interconnect_0:H0_s1_write -> H0:write_n
	wire  [31:0] mm_interconnect_0_h0_s1_writedata;                    // mm_interconnect_0:H0_s1_writedata -> H0:writedata
	wire         mm_interconnect_0_m1_s1_chipselect;                   // mm_interconnect_0:M1_s1_chipselect -> M1:chipselect
	wire  [31:0] mm_interconnect_0_m1_s1_readdata;                     // M1:readdata -> mm_interconnect_0:M1_s1_readdata
	wire   [1:0] mm_interconnect_0_m1_s1_address;                      // mm_interconnect_0:M1_s1_address -> M1:address
	wire         mm_interconnect_0_m1_s1_write;                        // mm_interconnect_0:M1_s1_write -> M1:write_n
	wire  [31:0] mm_interconnect_0_m1_s1_writedata;                    // mm_interconnect_0:M1_s1_writedata -> M1:writedata
	wire         mm_interconnect_0_m0_s1_chipselect;                   // mm_interconnect_0:M0_s1_chipselect -> M0:chipselect
	wire  [31:0] mm_interconnect_0_m0_s1_readdata;                     // M0:readdata -> mm_interconnect_0:M0_s1_readdata
	wire   [1:0] mm_interconnect_0_m0_s1_address;                      // mm_interconnect_0:M0_s1_address -> M0:address
	wire         mm_interconnect_0_m0_s1_write;                        // mm_interconnect_0:M0_s1_write -> M0:write_n
	wire  [31:0] mm_interconnect_0_m0_s1_writedata;                    // mm_interconnect_0:M0_s1_writedata -> M0:writedata
	wire         mm_interconnect_0_s1_s1_chipselect;                   // mm_interconnect_0:S1_s1_chipselect -> S1:chipselect
	wire  [31:0] mm_interconnect_0_s1_s1_readdata;                     // S1:readdata -> mm_interconnect_0:S1_s1_readdata
	wire   [1:0] mm_interconnect_0_s1_s1_address;                      // mm_interconnect_0:S1_s1_address -> S1:address
	wire         mm_interconnect_0_s1_s1_write;                        // mm_interconnect_0:S1_s1_write -> S1:write_n
	wire  [31:0] mm_interconnect_0_s1_s1_writedata;                    // mm_interconnect_0:S1_s1_writedata -> S1:writedata
	wire         mm_interconnect_0_s0_s1_chipselect;                   // mm_interconnect_0:S0_s1_chipselect -> S0:chipselect
	wire  [31:0] mm_interconnect_0_s0_s1_readdata;                     // S0:readdata -> mm_interconnect_0:S0_s1_readdata
	wire   [1:0] mm_interconnect_0_s0_s1_address;                      // mm_interconnect_0:S0_s1_address -> S0:address
	wire         mm_interconnect_0_s0_s1_write;                        // mm_interconnect_0:S0_s1_write -> S0:write_n
	wire  [31:0] mm_interconnect_0_s0_s1_writedata;                    // mm_interconnect_0:S0_s1_writedata -> S0:writedata
	wire         mm_interconnect_0_alarm_s1_chipselect;                // mm_interconnect_0:ALARM_s1_chipselect -> ALARM:chipselect
	wire  [31:0] mm_interconnect_0_alarm_s1_readdata;                  // ALARM:readdata -> mm_interconnect_0:ALARM_s1_readdata
	wire   [1:0] mm_interconnect_0_alarm_s1_address;                   // mm_interconnect_0:ALARM_s1_address -> ALARM:address
	wire         mm_interconnect_0_alarm_s1_write;                     // mm_interconnect_0:ALARM_s1_write -> ALARM:write_n
	wire  [31:0] mm_interconnect_0_alarm_s1_writedata;                 // mm_interconnect_0:ALARM_s1_writedata -> ALARM:writedata
	wire         mm_interconnect_0_btn_set_alarm_s1_chipselect;        // mm_interconnect_0:BTN_SET_ALARM_s1_chipselect -> BTN_SET_ALARM:chipselect
	wire  [31:0] mm_interconnect_0_btn_set_alarm_s1_readdata;          // BTN_SET_ALARM:readdata -> mm_interconnect_0:BTN_SET_ALARM_s1_readdata
	wire   [1:0] mm_interconnect_0_btn_set_alarm_s1_address;           // mm_interconnect_0:BTN_SET_ALARM_s1_address -> BTN_SET_ALARM:address
	wire         mm_interconnect_0_btn_set_alarm_s1_write;             // mm_interconnect_0:BTN_SET_ALARM_s1_write -> BTN_SET_ALARM:write_n
	wire  [31:0] mm_interconnect_0_btn_set_alarm_s1_writedata;         // mm_interconnect_0:BTN_SET_ALARM_s1_writedata -> BTN_SET_ALARM:writedata
	wire         mm_interconnect_0_btn_up_s1_chipselect;               // mm_interconnect_0:BTN_UP_s1_chipselect -> BTN_UP:chipselect
	wire  [31:0] mm_interconnect_0_btn_up_s1_readdata;                 // BTN_UP:readdata -> mm_interconnect_0:BTN_UP_s1_readdata
	wire   [1:0] mm_interconnect_0_btn_up_s1_address;                  // mm_interconnect_0:BTN_UP_s1_address -> BTN_UP:address
	wire         mm_interconnect_0_btn_up_s1_write;                    // mm_interconnect_0:BTN_UP_s1_write -> BTN_UP:write_n
	wire  [31:0] mm_interconnect_0_btn_up_s1_writedata;                // mm_interconnect_0:BTN_UP_s1_writedata -> BTN_UP:writedata
	wire         mm_interconnect_0_btn_down_s1_chipselect;             // mm_interconnect_0:BTN_DOWN_s1_chipselect -> BTN_DOWN:chipselect
	wire  [31:0] mm_interconnect_0_btn_down_s1_readdata;               // BTN_DOWN:readdata -> mm_interconnect_0:BTN_DOWN_s1_readdata
	wire   [1:0] mm_interconnect_0_btn_down_s1_address;                // mm_interconnect_0:BTN_DOWN_s1_address -> BTN_DOWN:address
	wire         mm_interconnect_0_btn_down_s1_write;                  // mm_interconnect_0:BTN_DOWN_s1_write -> BTN_DOWN:write_n
	wire  [31:0] mm_interconnect_0_btn_down_s1_writedata;              // mm_interconnect_0:BTN_DOWN_s1_writedata -> BTN_DOWN:writedata
	wire         mm_interconnect_0_btn_set_clock_s1_chipselect;        // mm_interconnect_0:BTN_SET_CLOCK_s1_chipselect -> BTN_SET_CLOCK:chipselect
	wire  [31:0] mm_interconnect_0_btn_set_clock_s1_readdata;          // BTN_SET_CLOCK:readdata -> mm_interconnect_0:BTN_SET_CLOCK_s1_readdata
	wire   [1:0] mm_interconnect_0_btn_set_clock_s1_address;           // mm_interconnect_0:BTN_SET_CLOCK_s1_address -> BTN_SET_CLOCK:address
	wire         mm_interconnect_0_btn_set_clock_s1_write;             // mm_interconnect_0:BTN_SET_CLOCK_s1_write -> BTN_SET_CLOCK:write_n
	wire  [31:0] mm_interconnect_0_btn_set_clock_s1_writedata;         // mm_interconnect_0:BTN_SET_CLOCK_s1_writedata -> BTN_SET_CLOCK:writedata
	wire         irq_mapper_receiver0_irq;                             // UART:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                             // BTN_SET_ALARM:irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                             // BTN_UP:irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                             // BTN_DOWN:irq -> irq_mapper:receiver3_irq
	wire         irq_mapper_receiver4_irq;                             // BTN_SET_CLOCK:irq -> irq_mapper:receiver4_irq
	wire  [31:0] cpu_irq_irq;                                          // irq_mapper:sender_irq -> CPU:irq
	wire         rst_controller_reset_out_reset;                       // rst_controller:reset_out -> [ALARM:reset_n, BTN_DOWN:reset_n, BTN_SET_ALARM:reset_n, BTN_SET_CLOCK:reset_n, BTN_UP:reset_n, CPU:reset_n, H0:reset_n, H1:reset_n, M0:reset_n, M1:reset_n, RAM:reset, S0:reset_n, S1:reset_n, UART:rst_n, irq_mapper:reset, mm_interconnect_0:CPU_reset_reset_bridge_in_reset_reset, rst_translator:in_reset]
	wire         rst_controller_reset_out_reset_req;                   // rst_controller:reset_req -> [CPU:reset_req, RAM:reset_req, rst_translator:reset_req_in]

	system_ALARM alarm (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_alarm_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_alarm_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_alarm_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_alarm_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_alarm_s1_readdata),   //                    .readdata
		.out_port   (alarm_export)                           // external_connection.export
	);

	system_BTN_DOWN btn_down (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_btn_down_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_btn_down_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_btn_down_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_btn_down_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_btn_down_s1_readdata),   //                    .readdata
		.in_port    (btn_down_export),                          // external_connection.export
		.irq        (irq_mapper_receiver3_irq)                  //                 irq.irq
	);

	system_BTN_DOWN btn_set_alarm (
		.clk        (clk_clk),                                       //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address    (mm_interconnect_0_btn_set_alarm_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_btn_set_alarm_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_btn_set_alarm_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_btn_set_alarm_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_btn_set_alarm_s1_readdata),   //                    .readdata
		.in_port    (btn_set_alarm_export),                          // external_connection.export
		.irq        (irq_mapper_receiver1_irq)                       //                 irq.irq
	);

	system_BTN_DOWN btn_set_clock (
		.clk        (clk_clk),                                       //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address    (mm_interconnect_0_btn_set_clock_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_btn_set_clock_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_btn_set_clock_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_btn_set_clock_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_btn_set_clock_s1_readdata),   //                    .readdata
		.in_port    (btn_set_clock_export),                          // external_connection.export
		.irq        (irq_mapper_receiver4_irq)                       //                 irq.irq
	);

	system_BTN_DOWN btn_up (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_btn_up_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_btn_up_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_btn_up_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_btn_up_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_btn_up_s1_readdata),   //                    .readdata
		.in_port    (btn_up_export),                          // external_connection.export
		.irq        (irq_mapper_receiver2_irq)                //                 irq.irq
	);

	system_CPU cpu (
		.clk                                 (clk_clk),                                           //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                   //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                //                          .reset_req
		.d_address                           (cpu_data_master_address),                           //               data_master.address
		.d_byteenable                        (cpu_data_master_byteenable),                        //                          .byteenable
		.d_read                              (cpu_data_master_read),                              //                          .read
		.d_readdata                          (cpu_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (cpu_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (cpu_data_master_write),                             //                          .write
		.d_writedata                         (cpu_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (cpu_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (cpu_instruction_master_address),                    //        instruction_master.address
		.i_read                              (cpu_instruction_master_read),                       //                          .read
		.i_readdata                          (cpu_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (cpu_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (cpu_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (),                                                  //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_cpu_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_cpu_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_cpu_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_cpu_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_cpu_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_cpu_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_cpu_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_cpu_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                   // custom_instruction_master.readra
	);

	system_H0 h0 (
		.clk        (clk_clk),                            //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),    //               reset.reset_n
		.address    (mm_interconnect_0_h0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_h0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_h0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_h0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_h0_s1_readdata),   //                    .readdata
		.out_port   (display_h0_export)                   // external_connection.export
	);

	system_H0 h1 (
		.clk        (clk_clk),                            //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),    //               reset.reset_n
		.address    (mm_interconnect_0_h1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_h1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_h1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_h1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_h1_s1_readdata),   //                    .readdata
		.out_port   (display_h1_export)                   // external_connection.export
	);

	system_H0 m0 (
		.clk        (clk_clk),                            //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),    //               reset.reset_n
		.address    (mm_interconnect_0_m0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_m0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_m0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_m0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_m0_s1_readdata),   //                    .readdata
		.out_port   (display_m0_export)                   // external_connection.export
	);

	system_H0 m1 (
		.clk        (clk_clk),                            //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),    //               reset.reset_n
		.address    (mm_interconnect_0_m1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_m1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_m1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_m1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_m1_s1_readdata),   //                    .readdata
		.out_port   (display_m1_export)                   // external_connection.export
	);

	system_RAM ram (
		.clk        (clk_clk),                             //   clk1.clk
		.address    (mm_interconnect_0_ram_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_ram_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_ram_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_ram_s1_write),      //       .write
		.readdata   (mm_interconnect_0_ram_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_ram_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_ram_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),      // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),  //       .reset_req
		.freeze     (1'b0)                                 // (terminated)
	);

	system_H0 s0 (
		.clk        (clk_clk),                            //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),    //               reset.reset_n
		.address    (mm_interconnect_0_s0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_s0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_s0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_s0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_s0_s1_readdata),   //                    .readdata
		.out_port   (display_s0_export)                   // external_connection.export
	);

	system_H0 s1 (
		.clk        (clk_clk),                            //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),    //               reset.reset_n
		.address    (mm_interconnect_0_s1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_s1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_s1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_s1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_s1_s1_readdata),   //                    .readdata
		.out_port   (display_s1_export)                   // external_connection.export
	);

	system_UART uart (
		.clk            (clk_clk),                                              //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                      //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                              //               irq.irq
	);

	system_mm_interconnect_0 mm_interconnect_0 (
		.CLK_clk_clk                           (clk_clk),                                              //                         CLK_clk.clk
		.CPU_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                       // CPU_reset_reset_bridge_in_reset.reset
		.CPU_data_master_address               (cpu_data_master_address),                              //                 CPU_data_master.address
		.CPU_data_master_waitrequest           (cpu_data_master_waitrequest),                          //                                .waitrequest
		.CPU_data_master_byteenable            (cpu_data_master_byteenable),                           //                                .byteenable
		.CPU_data_master_read                  (cpu_data_master_read),                                 //                                .read
		.CPU_data_master_readdata              (cpu_data_master_readdata),                             //                                .readdata
		.CPU_data_master_write                 (cpu_data_master_write),                                //                                .write
		.CPU_data_master_writedata             (cpu_data_master_writedata),                            //                                .writedata
		.CPU_data_master_debugaccess           (cpu_data_master_debugaccess),                          //                                .debugaccess
		.CPU_instruction_master_address        (cpu_instruction_master_address),                       //          CPU_instruction_master.address
		.CPU_instruction_master_waitrequest    (cpu_instruction_master_waitrequest),                   //                                .waitrequest
		.CPU_instruction_master_read           (cpu_instruction_master_read),                          //                                .read
		.CPU_instruction_master_readdata       (cpu_instruction_master_readdata),                      //                                .readdata
		.ALARM_s1_address                      (mm_interconnect_0_alarm_s1_address),                   //                        ALARM_s1.address
		.ALARM_s1_write                        (mm_interconnect_0_alarm_s1_write),                     //                                .write
		.ALARM_s1_readdata                     (mm_interconnect_0_alarm_s1_readdata),                  //                                .readdata
		.ALARM_s1_writedata                    (mm_interconnect_0_alarm_s1_writedata),                 //                                .writedata
		.ALARM_s1_chipselect                   (mm_interconnect_0_alarm_s1_chipselect),                //                                .chipselect
		.BTN_DOWN_s1_address                   (mm_interconnect_0_btn_down_s1_address),                //                     BTN_DOWN_s1.address
		.BTN_DOWN_s1_write                     (mm_interconnect_0_btn_down_s1_write),                  //                                .write
		.BTN_DOWN_s1_readdata                  (mm_interconnect_0_btn_down_s1_readdata),               //                                .readdata
		.BTN_DOWN_s1_writedata                 (mm_interconnect_0_btn_down_s1_writedata),              //                                .writedata
		.BTN_DOWN_s1_chipselect                (mm_interconnect_0_btn_down_s1_chipselect),             //                                .chipselect
		.BTN_SET_ALARM_s1_address              (mm_interconnect_0_btn_set_alarm_s1_address),           //                BTN_SET_ALARM_s1.address
		.BTN_SET_ALARM_s1_write                (mm_interconnect_0_btn_set_alarm_s1_write),             //                                .write
		.BTN_SET_ALARM_s1_readdata             (mm_interconnect_0_btn_set_alarm_s1_readdata),          //                                .readdata
		.BTN_SET_ALARM_s1_writedata            (mm_interconnect_0_btn_set_alarm_s1_writedata),         //                                .writedata
		.BTN_SET_ALARM_s1_chipselect           (mm_interconnect_0_btn_set_alarm_s1_chipselect),        //                                .chipselect
		.BTN_SET_CLOCK_s1_address              (mm_interconnect_0_btn_set_clock_s1_address),           //                BTN_SET_CLOCK_s1.address
		.BTN_SET_CLOCK_s1_write                (mm_interconnect_0_btn_set_clock_s1_write),             //                                .write
		.BTN_SET_CLOCK_s1_readdata             (mm_interconnect_0_btn_set_clock_s1_readdata),          //                                .readdata
		.BTN_SET_CLOCK_s1_writedata            (mm_interconnect_0_btn_set_clock_s1_writedata),         //                                .writedata
		.BTN_SET_CLOCK_s1_chipselect           (mm_interconnect_0_btn_set_clock_s1_chipselect),        //                                .chipselect
		.BTN_UP_s1_address                     (mm_interconnect_0_btn_up_s1_address),                  //                       BTN_UP_s1.address
		.BTN_UP_s1_write                       (mm_interconnect_0_btn_up_s1_write),                    //                                .write
		.BTN_UP_s1_readdata                    (mm_interconnect_0_btn_up_s1_readdata),                 //                                .readdata
		.BTN_UP_s1_writedata                   (mm_interconnect_0_btn_up_s1_writedata),                //                                .writedata
		.BTN_UP_s1_chipselect                  (mm_interconnect_0_btn_up_s1_chipselect),               //                                .chipselect
		.CPU_debug_mem_slave_address           (mm_interconnect_0_cpu_debug_mem_slave_address),        //             CPU_debug_mem_slave.address
		.CPU_debug_mem_slave_write             (mm_interconnect_0_cpu_debug_mem_slave_write),          //                                .write
		.CPU_debug_mem_slave_read              (mm_interconnect_0_cpu_debug_mem_slave_read),           //                                .read
		.CPU_debug_mem_slave_readdata          (mm_interconnect_0_cpu_debug_mem_slave_readdata),       //                                .readdata
		.CPU_debug_mem_slave_writedata         (mm_interconnect_0_cpu_debug_mem_slave_writedata),      //                                .writedata
		.CPU_debug_mem_slave_byteenable        (mm_interconnect_0_cpu_debug_mem_slave_byteenable),     //                                .byteenable
		.CPU_debug_mem_slave_waitrequest       (mm_interconnect_0_cpu_debug_mem_slave_waitrequest),    //                                .waitrequest
		.CPU_debug_mem_slave_debugaccess       (mm_interconnect_0_cpu_debug_mem_slave_debugaccess),    //                                .debugaccess
		.H0_s1_address                         (mm_interconnect_0_h0_s1_address),                      //                           H0_s1.address
		.H0_s1_write                           (mm_interconnect_0_h0_s1_write),                        //                                .write
		.H0_s1_readdata                        (mm_interconnect_0_h0_s1_readdata),                     //                                .readdata
		.H0_s1_writedata                       (mm_interconnect_0_h0_s1_writedata),                    //                                .writedata
		.H0_s1_chipselect                      (mm_interconnect_0_h0_s1_chipselect),                   //                                .chipselect
		.H1_s1_address                         (mm_interconnect_0_h1_s1_address),                      //                           H1_s1.address
		.H1_s1_write                           (mm_interconnect_0_h1_s1_write),                        //                                .write
		.H1_s1_readdata                        (mm_interconnect_0_h1_s1_readdata),                     //                                .readdata
		.H1_s1_writedata                       (mm_interconnect_0_h1_s1_writedata),                    //                                .writedata
		.H1_s1_chipselect                      (mm_interconnect_0_h1_s1_chipselect),                   //                                .chipselect
		.M0_s1_address                         (mm_interconnect_0_m0_s1_address),                      //                           M0_s1.address
		.M0_s1_write                           (mm_interconnect_0_m0_s1_write),                        //                                .write
		.M0_s1_readdata                        (mm_interconnect_0_m0_s1_readdata),                     //                                .readdata
		.M0_s1_writedata                       (mm_interconnect_0_m0_s1_writedata),                    //                                .writedata
		.M0_s1_chipselect                      (mm_interconnect_0_m0_s1_chipselect),                   //                                .chipselect
		.M1_s1_address                         (mm_interconnect_0_m1_s1_address),                      //                           M1_s1.address
		.M1_s1_write                           (mm_interconnect_0_m1_s1_write),                        //                                .write
		.M1_s1_readdata                        (mm_interconnect_0_m1_s1_readdata),                     //                                .readdata
		.M1_s1_writedata                       (mm_interconnect_0_m1_s1_writedata),                    //                                .writedata
		.M1_s1_chipselect                      (mm_interconnect_0_m1_s1_chipselect),                   //                                .chipselect
		.RAM_s1_address                        (mm_interconnect_0_ram_s1_address),                     //                          RAM_s1.address
		.RAM_s1_write                          (mm_interconnect_0_ram_s1_write),                       //                                .write
		.RAM_s1_readdata                       (mm_interconnect_0_ram_s1_readdata),                    //                                .readdata
		.RAM_s1_writedata                      (mm_interconnect_0_ram_s1_writedata),                   //                                .writedata
		.RAM_s1_byteenable                     (mm_interconnect_0_ram_s1_byteenable),                  //                                .byteenable
		.RAM_s1_chipselect                     (mm_interconnect_0_ram_s1_chipselect),                  //                                .chipselect
		.RAM_s1_clken                          (mm_interconnect_0_ram_s1_clken),                       //                                .clken
		.S0_s1_address                         (mm_interconnect_0_s0_s1_address),                      //                           S0_s1.address
		.S0_s1_write                           (mm_interconnect_0_s0_s1_write),                        //                                .write
		.S0_s1_readdata                        (mm_interconnect_0_s0_s1_readdata),                     //                                .readdata
		.S0_s1_writedata                       (mm_interconnect_0_s0_s1_writedata),                    //                                .writedata
		.S0_s1_chipselect                      (mm_interconnect_0_s0_s1_chipselect),                   //                                .chipselect
		.S1_s1_address                         (mm_interconnect_0_s1_s1_address),                      //                           S1_s1.address
		.S1_s1_write                           (mm_interconnect_0_s1_s1_write),                        //                                .write
		.S1_s1_readdata                        (mm_interconnect_0_s1_s1_readdata),                     //                                .readdata
		.S1_s1_writedata                       (mm_interconnect_0_s1_s1_writedata),                    //                                .writedata
		.S1_s1_chipselect                      (mm_interconnect_0_s1_s1_chipselect),                   //                                .chipselect
		.UART_avalon_jtag_slave_address        (mm_interconnect_0_uart_avalon_jtag_slave_address),     //          UART_avalon_jtag_slave.address
		.UART_avalon_jtag_slave_write          (mm_interconnect_0_uart_avalon_jtag_slave_write),       //                                .write
		.UART_avalon_jtag_slave_read           (mm_interconnect_0_uart_avalon_jtag_slave_read),        //                                .read
		.UART_avalon_jtag_slave_readdata       (mm_interconnect_0_uart_avalon_jtag_slave_readdata),    //                                .readdata
		.UART_avalon_jtag_slave_writedata      (mm_interconnect_0_uart_avalon_jtag_slave_writedata),   //                                .writedata
		.UART_avalon_jtag_slave_waitrequest    (mm_interconnect_0_uart_avalon_jtag_slave_waitrequest), //                                .waitrequest
		.UART_avalon_jtag_slave_chipselect     (mm_interconnect_0_uart_avalon_jtag_slave_chipselect)   //                                .chipselect
	);

	system_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),       // receiver4.irq
		.sender_irq    (cpu_irq_irq)                     //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
